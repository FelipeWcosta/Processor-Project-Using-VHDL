library verilog;
use verilog.vl_types.all;
entity processador_demonstracao_vlg_vec_tst is
end processador_demonstracao_vlg_vec_tst;
