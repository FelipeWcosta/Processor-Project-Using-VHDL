library verilog;
use verilog.vl_types.all;
entity ir_vlg_check_tst is
    port(
        IR_out          : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end ir_vlg_check_tst;
