library verilog;
use verilog.vl_types.all;
entity processador_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        rst_principal   : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end processador_vlg_sample_tst;
