library verilog;
use verilog.vl_types.all;
entity RF_Rp_vlg_vec_tst is
end RF_Rp_vlg_vec_tst;
