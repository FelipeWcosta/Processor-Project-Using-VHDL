library verilog;
use verilog.vl_types.all;
entity data_op_vlg_vec_tst is
end data_op_vlg_vec_tst;
