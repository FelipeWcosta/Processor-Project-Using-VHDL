library verilog;
use verilog.vl_types.all;
entity ir_vlg_vec_tst is
end ir_vlg_vec_tst;
