library verilog;
use verilog.vl_types.all;
entity data_i_vlg_vec_tst is
end data_i_vlg_vec_tst;
